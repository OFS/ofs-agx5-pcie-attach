// Copyright (C) 2021 Intel Corporation.
// SPDX-License-Identifier: MIT

//
// Description
//-----------------------------------------------------------------------------
//
// This package defines the global parameters of FIM
//
//----------------------------------------------------------------------------

`ifndef __OFS_FIM_CFG_PKG_SV__
`define __OFS_FIM_CFG_PKG_SV__

// IP configuration database, generated by OFS script ofs_ip_cfg_db.tcl after
// IP generation.
`include "ofs_ip_cfg_db.vh"

package ofs_fim_cfg_pkg;

localparam real MAIN_CLK_MHZ = sys_pll_pkg::clock_name_to_actual_mhz("clk_sys");

//*****************
// PCIe host parameters
//*****************
localparam PCIE_LANES = `OFS_FIM_IP_CFG_PCIE_SS_TOTAL_NUM_LANES;

localparam NUM_PCIE_HOST      = 1;
localparam PCIE_HOST_WIDTH    = $clog2(NUM_PCIE_HOST);

// Native width of the AXI-S TLP stream from the PCIe IP
localparam PCIE_IP_TDATA_WIDTH = `OFS_FIM_IP_CFG_PCIE_SS_DWIDTH_BYTE * 8;
// Width of the OFS internal TLP stream. May be transformed to a value
// different from the IP itself. OFS requires a PCIe bus at least wide enough
// to hold a complete TLP header.
localparam PCIE_TDATA_WIDTH  = (PCIE_IP_TDATA_WIDTH >= 256) ? PCIE_IP_TDATA_WIDTH : 256;
localparam PCIE_TUSER_WIDTH  = 10;
localparam PCIE_LITE_CSR_WIDTH = 20;

localparam PCIE_RP_MAX_TAGS   = (1<<10);
localparam PCIE_RP_TAG_WIDTH  = $clog2(PCIE_RP_MAX_TAGS);

localparam MAX_PAYLOAD_SIZE   = 128; // DW
localparam MAX_RD_REQ_SIZE    = 128; // DW

`ifdef OFS_FIM_IP_CFG_PCIE_SS_FUNC_MODE_IS_DM
  localparam PCIE_DM_ENCODING_EN = 1;
`else
  localparam PCIE_DM_ENCODING_EN = 0;
`endif

`ifdef OFS_FIM_IP_CFG_PCIE_SS_HAS_CPL_REORDER
  localparam PCIE_CPL_REORDER_EN = 1;
`else
  localparam PCIE_CPL_REORDER_EN = 0;
`endif

//*****************
// MMIO parameters
//*****************
localparam PORTS              = 1;
localparam MMIO_TID_WIDTH     = PCIE_HOST_WIDTH + PCIE_RP_TAG_WIDTH; // Matches PCIe TLP tag width 
localparam MMIO_DATA_WIDTH    = 64;
// PF0 bar 0 addr width 1MB, VF under this PF has same address width
localparam MMIO_ADDR_WIDTH    = `OFS_FIM_IP_CFG_PCIE_SS_PF0_BAR0_ADDR_WIDTH;
// PF0 BAR0 VF address width
`ifdef OFS_FIM_IP_CFG_PCIE_SS_PF0_VF_BAR0_ADDR_WIDTH
  localparam MMIO_ADDR_WIDTH_PG = `OFS_FIM_IP_CFG_PCIE_SS_PF0_VF_BAR0_ADDR_WIDTH;
`else
  localparam MMIO_ADDR_WIDTH_PG = MMIO_ADDR_WIDTH;  // Pick a default
`endif 
// non PF0 bar 0 (often 4KB)
`ifdef OFS_FIM_IP_CFG_PCIE_SS_PF1_BAR0_ADDR_WIDTH
  localparam NONPF0_MMIO_ADDR_WIDTH = `OFS_FIM_IP_CFG_PCIE_SS_PF1_BAR0_ADDR_WIDTH;
`else
  localparam NONPF0_MMIO_ADDR_WIDTH = 12;  // Pick a default
`endif

`ifdef NUM_AFUS
localparam   NUM_AFUS    = 2;
`else
localparam   NUM_AFUS    = 1;
`endif
localparam LNUM_AFUS = NUM_AFUS>1?$clog2(NUM_AFUS):1'h1;


// MSIX

// Number of interrupts is encoded per-PF/VF from the PCIe IP as a vector
localparam int MSIX_PF_TABLE_SIZE[8] = '{ `OFS_FIM_IP_CFG_PCIE_SS_MSIX_PF_TABLE_SIZE_VEC };
localparam int MSIX_VF_TABLE_SIZE[8] = '{ `OFS_FIM_IP_CFG_PCIE_SS_MSIX_VF_TABLE_SIZE_VEC };

// OFS expects each function to have the same MSI-X configuration.
// Try VF0. Failing that, use PF0.
localparam NUM_AFU_INTERRUPTS = MSIX_VF_TABLE_SIZE[0] ? MSIX_VF_TABLE_SIZE[0] : MSIX_PF_TABLE_SIZE[0];
localparam L_NUM_AFU_INTERRUPTS = $clog2(NUM_AFU_INTERRUPTS);

endpackage

`endif // __OFS_FIM_CFG_PKG_SV__
